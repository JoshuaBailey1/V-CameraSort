module camsort_modules

pub fn do_nothing()
{
	
}